--#############################################################################
-- institute: BTU
--
-- author: Keyvan Shahin
--
-- date: Sep, 15, 2021
--
--#############################################################################

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package parameters is
	
	--WRD related
	constant cIWGlobal		: integer := 16; --Input Integer part Width
	constant cFWGlobal		: integer := 16; --Input Integer part Width
	--constant cAddSubSel		: boolean := true; --true for add, false for sub
	
	subtype tIntWidth	is integer range 0 to cIWGlobal;
	subtype tFloatWidth	is integer range 0 to cFWGlobal;
	
	--FIR Related
	constant cNumberOfTaps : integer := 51;	-- number of FIR taps

	type	tIntWidthArray is array (natural range <>) of tIntWidth;
	type	tFloatWidthArray is array (natural range <>) of tFloatWidth;
	
	subtype	tDataPath	is signed (cIWGlobal+cFWGlobal-1 downto 0);
	type	tDataPathArray	is array (natural range <>) of tDataPath; --Delay Line Type
	constant cCoeff	: tDataPathArray (cNumberOfTaps-1 downto 0);
end package parameters;

package body parameters is 
	--FIR Coefficients
	constant cCoeff	: tDataPathArray (cNumberOfTaps-1 downto 0) := 
	(
	"00000000000000010000000000000000",
	"00000000000000010000000000000000",
	"00000000000000010000000000000000",
	"00000000000000010000000000000000",
	"00000000000000010000000000000000",
	"00000000000000010000000000000000",
	"00000000000000010000000000000000",
	"00000000000000010000000000000000",
	"00000000000000010000000000000000",
	"00000000000000010000000000000000",
	"00000000000000010000000000000000",
	"00000000000000010000000000000000",
	"00000000000000010000000000000000",
	"00000000000000010000000000000000",
	"00000000000000010000000000000000",
	"00000000000000010000000000000000",
	"00000000000000010000000000000000",
	"00000000000000010000000000000000",
	"00000000000000010000000000000000",
	"00000000000000010000000000000000",
	"00000000000000010000000000000000",
	"00000000000000010000000000000000",
	"00000000000000010000000000000000",
	"00000000000000010000000000000000",
	"00000000000000010000000000000000",
	"00000000000000010000000000000000",
	"00000000000000010000000000000000",
	"00000000000000010000000000000000",
	"00000000000000010000000000000000",
	"00000000000000010000000000000000",
	"00000000000000010000000000000000",
	"00000000000000010000000000000000",
	"00000000000000010000000000000000",
	"00000000000000010000000000000000",
	"00000000000000010000000000000000",
	"00000000000000010000000000000000",
	"00000000000000010000000000000000",
	"00000000000000010000000000000000",
	"00000000000000010000000000000000",
	"00000000000000010000000000000000",
	"00000000000000010000000000000000",
	"00000000000000010000000000000000",
	"00000000000000010000000000000000",
	"00000000000000010000000000000000",
	"00000000000000010000000000000000",
	"00000000000000010000000000000000",
	"00000000000000010000000000000000",
	"00000000000000010000000000000000",
	"00000000000000010000000000000000",
	"00000000000000010000000000000000",
	"00000000000000010000000000000000"
	);
end package body parameters; 
